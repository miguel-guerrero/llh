module Const(z);

parameter W=1;
parameter VAL=0;

output [W-1:0] z;

assign z = VAL;

endmodule
